library IEEE;
use IEEE.STD_LOGIC_1164.all;

ENTITY MUX2_4W_with_select_when IS 
PORT(X:IN STD_LOGIC_VECTOR(1 downto 0);
		D0,D1,D2,D3:IN STD_LOGIC;
		LED_COM:out std_logic;
		Y:OUT STD_LOGIC);
END MUX2_4W_with_select_when;

ARCHITECTURE mux2to4w OF MUX2_4W_with_select_when IS
BEGIN 
	LED_COM<='1';
	With X select
	 Y<=D0 when "00",
		D1 when "01",
		D2 when "10",
		D3 when others;
END mux2to4w;